module and_gate (
    input wire a,    // First input
    input wire b,    // Second input
    output wire y    // Output
);

    assign y = a & b; // AND operation

endmodule
